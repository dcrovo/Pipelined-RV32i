--PONTIFICIA_UNIVERSIDAD_JAVERIANA-- 
--VHDL DE ALU DE RVI32--
--DISEÑADOR: DANIEL_FAJARDO--
--6/10/2020--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

--En esta seccion se colocan las senales de entrada y salidas basandonos en el diagrama en bloques.
entity ALU32 is
       port( Salida_ALU1 : out STD_LOGIC_VECTOR(31 downto 0);
				 Salida_ALU2 : out STD_LOGIC;
				 ALU_Control : in STD_LOGIC_VECTOR(2 downto 0);
				 ALU_Control2 : in STD_LOGIC_VECTOR(3 downto 0);--En el caso de que no sea una instruccion tipo R se debe realiar una extension de signo.
		       Salida_IRMux: in STD_LOGIC_VECTOR(31 downto 0);--Salida_IRMux---->A
				 Salida_BR_OUT1 : in STD_LOGIC_VECTOR(31 downto 0);--Salida_BR_OUT2------>B
				 --------PRUEBAS--
				 --mayor: out STD_LOGIC;
				 --menor: out STD_LOGIC;
				 --igual: out STD_LOGIC;
				 --noigual: out STD_LOGIC;
				 --restasalida: out STD_LOGIC_VECTOR(31 downto 0);
				 --twocomple: out STD_LOGIC_VECTOR(31 downto 0);
				 --onecomple: out STD_LOGIC_VECTOR(31 downto 0);
				 ---------------------------------------------
				 
		       Exce_ALU :in STD_LOGIC);
end ALU32;

architecture ALU32Arch of ALU32 is
signal AlmacenamientoA: std_logic_vector(31 downto 0);
signal AlmacenamientoB: std_logic_vector(31 downto 0);
signal AlmacenamientoBN: std_logic_vector(31 downto 0);
signal complemento1: std_logic_vector(31 downto 0);
signal complemento2: std_logic_vector(31 downto 0);
signal Resultado1: std_logic_vector(31 downto 0);
signal Resultado2: std_logic_vector(31 downto 0);
signal Resultado3: std_logic_vector(31 downto 0);
signal Resultado4: std_logic_vector(31 downto 0);
signal Resultado5: std_logic_vector(31 downto 0);
signal Resultado6: std_logic_vector(31 downto 0);
signal Resultado7: std_logic_vector(31 downto 0);
signal Salida1: std_logic_vector(31 downto 0);
signal Salida2: std_logic_vector(31 downto 0);
signal Salida3: std_logic_vector(31 downto 0);
signal Salida4: std_logic_vector(31 downto 0);
signal Salida5: std_logic_vector(31 downto 0);
signal Salida6 :std_logic_vector(31 downto 0);
signal Salida7 :std_logic_vector(31 downto 0);
signal Acarreo :std_logic_vector(31 downto 0);

 

signal OpcodeSuma,OpCodeResta,OpcodeOr,OpcodeAnd,OpcodeXor,Equal_Than,Less_Than,Larger_Than,OpcodeRotate,OpcodeShift,Not_Equal_Than: std_logic;

signal Carry0, Carry1,Carry2,Carry3,Carry4,Carry5,Carry6,Carry7,Carry8,Carry9,Carry10,Carry11,Carry12,Carry13,Carry14,Carry15,Carry16,Carry17,Carry18,
Carry19, Carry20,Carry21,Carry22,Carry23,Carry24,Carry25,Carry26,Carry27,Carry28,Carry29,Carry30,CarryZ0, CarryZ1,CarryZ2,CarryZ3,CarryZ4,CarryZ5,CarryZ6,CarryZ7,CarryZ8,CarryZ9,CarryZ10,CarryZ11,CarryZ12,CarryZ13,CarryZ14,CarryZ15,CarryZ16,CarryZ17,CarryZ18,
CarryZ19, CarryZ20,CarryZ21,CarryZ22,CarryZ23,CarryZ24,CarryZ25,CarryZ26,CarryZ27,CarryZ28,CarryZ29,CarryZ30,CarryX0, CarryX1,CarryX2,CarryX3,CarryX4,CarryX5,CarryX6,CarryX7,CarryX8,CarryX9,CarryX10,CarryX11,CarryX12,CarryX13,CarryX14,CarryX15,CarryX16,CarryX17,CarryX18,
CarryX19, CarryX20,CarryX21,CarryX22,CarryX23,CarryX24,CarryX25,CarryX26,CarryX27,CarryX28,CarryX29,CarryX30: std_logic; --Señales de 1 bit

signal AlmacI :std_logic;
 begin
 
 
 Acarreo(0)<='1';
 Acarreo(1)<='0';
 Acarreo(2)<='0';
 Acarreo(3)<='0';
 Acarreo(4)<='0';
 Acarreo(5)<='0';
 Acarreo(6)<='0';
 Acarreo(7)<='0';
 Acarreo(8)<='0';
 Acarreo(9)<='0';
 Acarreo(10)<='0';
 Acarreo(11)<='0';
 Acarreo(12)<='0';
 Acarreo(13)<='0';
 Acarreo(14)<='0';
 Acarreo(15)<='0';
 Acarreo(16)<='0';		 
 Acarreo(17)<='0';
 Acarreo(18)<='0';
 Acarreo(19)<='0';
 Acarreo(20)<='0';
 Acarreo(21)<='0';
 Acarreo(22)<='0';
 Acarreo(23)<='0';
 Acarreo(24)<='0';
 Acarreo(25)<='0';		 
 Acarreo(26)<='0';
 Acarreo(27)<='0';
 Acarreo(28)<='0';
 Acarreo(29)<='0';
 Acarreo(30)<='0';
 Acarreo(31)<='0';

-----------La senal Exce_ALU habilita el paso de Data--------
AlmacenamientoA(0)  <= Salida_IRMux(0) and  Exce_ALU;  
AlmacenamientoA(1)  <= Salida_IRMux(1) and Exce_ALU;    
AlmacenamientoA(2)  <= Salida_IRMux(2) and Exce_ALU;    
AlmacenamientoA(3)  <= Salida_IRMux(3) and Exce_ALU;    
AlmacenamientoA(4)  <= Salida_IRMux(4) and Exce_ALU;    
AlmacenamientoA(5)  <= Salida_IRMux(5) and Exce_ALU;    
AlmacenamientoA(6)  <= Salida_IRMux(6) and Exce_ALU;    
AlmacenamientoA(7)  <= Salida_IRMux(7) and Exce_ALU;    
AlmacenamientoA(8)  <= Salida_IRMux(8) and Exce_ALU;    
AlmacenamientoA(9)  <= Salida_IRMux(9) and Exce_ALU;    
AlmacenamientoA(10)  <= Salida_IRMux(10) and Exce_ALU;    
AlmacenamientoA(11)  <= Salida_IRMux(11) and Exce_ALU;    
AlmacenamientoA(12)  <= Salida_IRMux(12) and Exce_ALU;    
AlmacenamientoA(13)  <= Salida_IRMux(13) and Exce_ALU;    
AlmacenamientoA(14)  <= Salida_IRMux(14) and Exce_ALU;    
AlmacenamientoA(15)  <= Salida_IRMux(15) and Exce_ALU;    
AlmacenamientoA(16)  <= Salida_IRMux(16) and Exce_ALU;    
AlmacenamientoA(17)  <= Salida_IRMux(17) and Exce_ALU;   
AlmacenamientoA(18)  <= Salida_IRMux(18) and Exce_ALU;    
AlmacenamientoA(19)  <= Salida_IRMux(19) and Exce_ALU;    
AlmacenamientoA(20)  <= Salida_IRMux(20) and Exce_ALU;    
AlmacenamientoA(21)  <= Salida_IRMux(21) and Exce_ALU;    
AlmacenamientoA(22)  <= Salida_IRMux(22) and Exce_ALU;    
AlmacenamientoA(23)  <= Salida_IRMux(23) and Exce_ALU;    
AlmacenamientoA(24)  <= Salida_IRMux(24) and Exce_ALU;    
AlmacenamientoA(25)  <= Salida_IRMux(25) and Exce_ALU;    
AlmacenamientoA(26)  <= Salida_IRMux(26) and Exce_ALU;    
AlmacenamientoA(27)  <= Salida_IRMux(27) and Exce_ALU;    
AlmacenamientoA(28)  <= Salida_IRMux(28) and Exce_ALU;    
AlmacenamientoA(29)  <= Salida_IRMux(29) and Exce_ALU;    
AlmacenamientoA(30)  <= Salida_IRMux(30) and Exce_ALU;    
AlmacenamientoA(31)  <= Salida_IRMux(31) and Exce_ALU;

AlmacenamientoB(0)  <= Salida_BR_OUT1(0) and  Exce_ALU;  
AlmacenamientoB(1)  <= Salida_BR_OUT1(1) and Exce_ALU;    
AlmacenamientoB(2)  <= Salida_BR_OUT1(2) and Exce_ALU;    
AlmacenamientoB(3)  <= Salida_BR_OUT1(3) and Exce_ALU;    
AlmacenamientoB(4)  <= Salida_BR_OUT1(4) and Exce_ALU;    
AlmacenamientoB(5)  <= Salida_BR_OUT1(5) and Exce_ALU;    
AlmacenamientoB(6)  <= Salida_BR_OUT1(6) and Exce_ALU;    
AlmacenamientoB(7)  <= Salida_BR_OUT1(7) and Exce_ALU;    
AlmacenamientoB(8)  <= Salida_BR_OUT1(8) and Exce_ALU;    
AlmacenamientoB(9)  <= Salida_BR_OUT1(9) and Exce_ALU;    
AlmacenamientoB(10)  <= Salida_BR_OUT1(10) and Exce_ALU;    
AlmacenamientoB(11)  <= Salida_BR_OUT1(11) and Exce_ALU;    
AlmacenamientoB(12)  <= Salida_BR_OUT1(12) and Exce_ALU;    
AlmacenamientoB(13)  <= Salida_BR_OUT1(13) and Exce_ALU;    
AlmacenamientoB(14)  <= Salida_BR_OUT1(14) and Exce_ALU;    
AlmacenamientoB(15)  <= Salida_BR_OUT1(15) and Exce_ALU;    
AlmacenamientoB(16)  <= Salida_BR_OUT1(16) and Exce_ALU;    
AlmacenamientoB(17)  <= Salida_BR_OUT1(17) and Exce_ALU;   
AlmacenamientoB(18)  <= Salida_BR_OUT1(18) and Exce_ALU;    
AlmacenamientoB(19)  <= Salida_BR_OUT1(19) and Exce_ALU;    
AlmacenamientoB(20)  <= Salida_BR_OUT1(20) and Exce_ALU;    
AlmacenamientoB(21)  <= Salida_BR_OUT1(21) and Exce_ALU;    
AlmacenamientoB(22)  <= Salida_BR_OUT1(22) and Exce_ALU;    
AlmacenamientoB(23)  <= Salida_BR_OUT1(23) and Exce_ALU;    
AlmacenamientoB(24)  <= Salida_BR_OUT1(24) and Exce_ALU;    
AlmacenamientoB(25)  <= Salida_BR_OUT1(25) and Exce_ALU;    
AlmacenamientoB(26)  <= Salida_BR_OUT1(26) and Exce_ALU;    
AlmacenamientoB(27)  <= Salida_BR_OUT1(27) and Exce_ALU;    
AlmacenamientoB(28)  <= Salida_BR_OUT1(28) and Exce_ALU;    
AlmacenamientoB(29)  <= Salida_BR_OUT1(29) and Exce_ALU;    
AlmacenamientoB(30)  <= Salida_BR_OUT1(30) and Exce_ALU;    
AlmacenamientoB(31)  <= Salida_BR_OUT1(31) and Exce_ALU;

----------------Se niega las entradas para la resta------
AlmacenamientoBN(0)  <=not AlmacenamientoB(0) ;
AlmacenamientoBN(1)  <= not AlmacenamientoB(1);
AlmacenamientoBN(2)  <= not AlmacenamientoB(2);
AlmacenamientoBN(3)  <= not AlmacenamientoB(3);
AlmacenamientoBN(4)  <= not AlmacenamientoB(4);    
AlmacenamientoBN(5)  <= not AlmacenamientoB(5);
AlmacenamientoBN(6)  <= not AlmacenamientoB(6);
AlmacenamientoBN(7)  <= not AlmacenamientoB(7);
AlmacenamientoBN(8)  <= not AlmacenamientoB(8);
AlmacenamientoBN(9)  <= not AlmacenamientoB(9);
AlmacenamientoBN(10)  <= not AlmacenamientoB(10);
AlmacenamientoBN(11)  <= not AlmacenamientoB(11);
AlmacenamientoBN(12)  <= not AlmacenamientoB(12);
AlmacenamientoBN(13)  <= not AlmacenamientoB(13);
AlmacenamientoBN(14)  <= not AlmacenamientoB(14);
AlmacenamientoBN(15)  <= not AlmacenamientoB(15);
AlmacenamientoBN(16)  <= not AlmacenamientoB(16);
AlmacenamientoBN(17)  <= not AlmacenamientoB(17);
AlmacenamientoBN(18)  <= not AlmacenamientoB(18);
AlmacenamientoBN(19)  <= not AlmacenamientoB(19);
AlmacenamientoBN(20)  <= not AlmacenamientoB(20);
AlmacenamientoBN(21)  <= not AlmacenamientoB(21);
AlmacenamientoBN(22)  <= not AlmacenamientoB(22);
AlmacenamientoBN(23)  <= not AlmacenamientoB(23);    
AlmacenamientoBN(24)  <= not AlmacenamientoB(24);
AlmacenamientoBN(25)  <= not AlmacenamientoB(25);
AlmacenamientoBN(26)  <= not AlmacenamientoB(26);     
AlmacenamientoBN(27)  <= not AlmacenamientoB(27);    
AlmacenamientoBN(28)  <= not AlmacenamientoB(28);    
AlmacenamientoBN(29)  <= not AlmacenamientoB(29);
AlmacenamientoBN(30)  <= not AlmacenamientoB(30);    
AlmacenamientoBN(31)  <= not AlmacenamientoB(31);

 AlmacI<='1';
 
--------------ALU------------------------

----------SUM-------
Resultado1(0) <= ((AlmacenamientoA(0) and (AlmacenamientoB(0)xnor not AlmacI)) or (not AlmacenamientoA(0) and (AlmacenamientoB(0) xor not AlmacI))); 
Carry0 <= (AlmacenamientoA(0) and (AlmacenamientoB(0)));  

Resultado1(1) <= (AlmacenamientoA(1) and (AlmacenamientoB(1) xnor Carry0)) or (not AlmacenamientoA(1) and (AlmacenamientoB(1) xor Carry0)); 
Carry1 <= (AlmacenamientoA(1) and (AlmacenamientoB(1) xor Carry0)) or (AlmacenamientoB(1) and Carry0); 

Resultado1(2) <= (AlmacenamientoA(2)and (AlmacenamientoB(2)xnor Carry1)) or (not AlmacenamientoA(2)and (AlmacenamientoB(2)xor Carry1)); 
Carry2 <= (AlmacenamientoA(2)and (AlmacenamientoB(2)xor Carry1)) or (AlmacenamientoB(2)and Carry1); 

Resultado1(3) <= (AlmacenamientoA(3)and (AlmacenamientoB(3)xnor Carry2)) or (not AlmacenamientoA(3)and  (AlmacenamientoB(3)xor Carry2)); 
Carry3 <= (AlmacenamientoA(3)and (AlmacenamientoB(3)xor Carry2)) or (AlmacenamientoB(3)and Carry2); 

Resultado1(4) <= (AlmacenamientoA(4)and (AlmacenamientoB(4)xnor Carry3)) or (not AlmacenamientoA(4)and (AlmacenamientoB(4)xor Carry3)); 
Carry4 <= (AlmacenamientoA(4)and (AlmacenamientoB(4)xor Carry3)) or (AlmacenamientoB(4)and Carry3); 

Resultado1(5) <= (AlmacenamientoA(5) and (AlmacenamientoB(5) xnor Carry4)) or (not AlmacenamientoA(5) and (AlmacenamientoB(5) xor Carry4)); 
Carry5 <= (AlmacenamientoA(5) and (AlmacenamientoB(5) xor Carry4)) or (AlmacenamientoB(5) and Carry4); 

Resultado1(6) <= (AlmacenamientoA(6) and (AlmacenamientoB(6) xnor Carry5)) or (not AlmacenamientoA(6) and (AlmacenamientoB(6) xor Carry5)); 
Carry6 <= (AlmacenamientoA(6) and (AlmacenamientoB(6) xor Carry5)) or (AlmacenamientoB(6) and Carry5); 

Resultado1(7) <= (AlmacenamientoA(7) and (AlmacenamientoB(7) xnor Carry6)) or (not AlmacenamientoA(7) and (AlmacenamientoB(7) xor Carry6)); 
Carry7 <= (AlmacenamientoA(7) and (AlmacenamientoB(7) xor Carry6)) or (AlmacenamientoB(7) and Carry6); 

Resultado1(8) <= (AlmacenamientoA(8) and (AlmacenamientoB(8) xnor Carry7)) or (not AlmacenamientoA(8) and (AlmacenamientoB(8) xor Carry7)); 
Carry8 <= (AlmacenamientoA(8) and (AlmacenamientoB(8) xor Carry7)) or (AlmacenamientoB(8) and Carry7); 

Resultado1(9) <= (AlmacenamientoA(9) and (AlmacenamientoB(9) xnor Carry8)) or (not AlmacenamientoA(9) and (AlmacenamientoB(9) xor Carry8));
Carry9 <= (AlmacenamientoA(9) and (AlmacenamientoB(9) xor Carry8)) or (AlmacenamientoB(9) and Carry8); 

Resultado1(10) <= (AlmacenamientoA(10) and (AlmacenamientoB(10) xnor Carry9)) or (not AlmacenamientoA(10) and (AlmacenamientoB(10) xor Carry9)); 
Carry10 <= (AlmacenamientoA(10) and (AlmacenamientoB(10) xor Carry9)) or (AlmacenamientoB(10) and Carry9); 

Resultado1(11) <= (AlmacenamientoA(11) and (AlmacenamientoB(11) xnor Carry10)) or (not AlmacenamientoA(11) and (AlmacenamientoB(11) xor Carry10)); 
Carry11 <= (AlmacenamientoA(11) and (AlmacenamientoB(11) xor Carry10)) or (AlmacenamientoB(11) and Carry10); 

Resultado1(12) <= (AlmacenamientoA(12) and (AlmacenamientoB(12) xnor Carry11)) or (not AlmacenamientoA(12) and (AlmacenamientoB(12) xor Carry11)); 
Carry12 <= (AlmacenamientoA(12) and (AlmacenamientoB(12) xor Carry11)) or (AlmacenamientoB(12) and Carry11); 

Resultado1(13) <= (AlmacenamientoA(13) and (AlmacenamientoB(13) xnor Carry12)) or (not AlmacenamientoA(13) and (AlmacenamientoB(13) xor Carry12)); 
Carry13 <= (AlmacenamientoA(13) and (AlmacenamientoB(13) xor Carry12)) or (AlmacenamientoB(13) and Carry12); 

Resultado1(14) <= (AlmacenamientoA(14) and (AlmacenamientoB(14) xnor Carry13)) or (not AlmacenamientoA(14) and (AlmacenamientoB(14) xor Carry13)); 
Carry14 <= (AlmacenamientoA(14) and (AlmacenamientoB(14) xor Carry13)) or (AlmacenamientoB(14) and Carry13); 
 
Resultado1(15) <= (AlmacenamientoA(15) and (AlmacenamientoB(15) xnor Carry14)) or (not AlmacenamientoA(15) and (AlmacenamientoB(15) xor Carry14)); 
Carry15 <= (AlmacenamientoA(15) and (AlmacenamientoB(15) xor Carry14)) or (AlmacenamientoB(15) and Carry14); 

Resultado1(16) <= (AlmacenamientoA(16) and (AlmacenamientoB(16) xnor Carry15)) or (not AlmacenamientoA(16) and (AlmacenamientoB(16) xor Carry15)); 
Carry16 <= (AlmacenamientoA(16) and (AlmacenamientoB(16) xor Carry15)) or (AlmacenamientoB(16) and Carry15); 

Resultado1(17) <= (AlmacenamientoA(17)and (AlmacenamientoB(17)xnor Carry16)) or (not AlmacenamientoA(17)and (AlmacenamientoB(17)xor Carry16)); 
Carry17 <= (AlmacenamientoA(17)and (AlmacenamientoB(17)xor Carry16)) or (AlmacenamientoB(17)and Carry16); 

Resultado1(18) <= (AlmacenamientoA(18)and (AlmacenamientoB(18)xnor Carry17)) or (not AlmacenamientoA(18)and  (AlmacenamientoB(18)xor Carry17)); 
Carry18<= (AlmacenamientoA(18)and (AlmacenamientoB(18)xor Carry17)) or (AlmacenamientoB(18)and Carry17); 

Resultado1(19) <= (AlmacenamientoA(19)and (AlmacenamientoB(19)xnor Carry18)) or (not AlmacenamientoA(19)and (AlmacenamientoB(19)xor Carry18)); 
Carry19 <= (AlmacenamientoA(19)and (AlmacenamientoB(19)xor Carry18)) or (AlmacenamientoB(19)and Carry18); 

Resultado1(20) <= (AlmacenamientoA(20) and (AlmacenamientoB(20) xnor Carry19)) or (not AlmacenamientoA(20) and (AlmacenamientoB(20) xor Carry19)); 
Carry20 <= (AlmacenamientoA(20) and (AlmacenamientoB(20) xor Carry19)) or (AlmacenamientoB(20) and Carry19); 

Resultado1(21) <= (AlmacenamientoA(21) and (AlmacenamientoB(21) xnor Carry20)) or (not AlmacenamientoA(21) and (AlmacenamientoB(21) xor Carry20)); 
Carry21 <= (AlmacenamientoA(21) and (AlmacenamientoB(21) xor Carry20)) or (AlmacenamientoB(21) and Carry20); 

Resultado1(22) <= (AlmacenamientoA(22) and (AlmacenamientoB(22) xnor Carry21)) or (not AlmacenamientoA(22) and (AlmacenamientoB(22) xor Carry21)); 
Carry22 <= (AlmacenamientoA(22) and (AlmacenamientoB(22) xor Carry21)) or (AlmacenamientoB(22) and Carry21); 

Resultado1(23) <= (AlmacenamientoA(23) and (AlmacenamientoB(23) xnor Carry22)) or (not AlmacenamientoA(23) and (AlmacenamientoB(23) xor Carry22)); 
Carry23 <= (AlmacenamientoA(23) and (AlmacenamientoB(23) xor Carry22)) or (AlmacenamientoB(23) and Carry22); 
 
Resultado1(24) <= (AlmacenamientoA(24) and (AlmacenamientoB(24) xnor Carry23)) or (not AlmacenamientoA(24) and (AlmacenamientoB(24) xor Carry23)); 
Carry24 <= (AlmacenamientoA(24) and (AlmacenamientoB(24) xor Carry23)) or (AlmacenamientoB(24) and Carry23); 

Resultado1(25) <= (AlmacenamientoA(25) and (AlmacenamientoB(25) xnor Carry24)) or (not AlmacenamientoA(25) and (AlmacenamientoB(25) xor Carry24)); 
Carry25 <= (AlmacenamientoA(25) and (AlmacenamientoB(25) xor Carry24)) or (AlmacenamientoB(25) and Carry24); 

Resultado1(26) <= (AlmacenamientoA(26) and (AlmacenamientoB(26) xnor Carry25)) or (not AlmacenamientoA(26) and (AlmacenamientoB(26) xor Carry25)); 
Carry26 <= (AlmacenamientoA(26) and (AlmacenamientoB(26) xor Carry25)) or (AlmacenamientoB(26) and Carry25); 

Resultado1(27) <= (AlmacenamientoA(27) and (AlmacenamientoB(27) xnor Carry26)) or (not AlmacenamientoA(27) and (AlmacenamientoB(27) xor Carry26)); 
Carry27 <= (AlmacenamientoA(27) and (AlmacenamientoB(27) xor Carry26)) or (AlmacenamientoB(27) and Carry26); 

Resultado1(28) <= (AlmacenamientoA(28) and (AlmacenamientoB(28) xnor Carry27)) or (not AlmacenamientoA(28) and (AlmacenamientoB(28) xor Carry27)); 
Carry28 <= (AlmacenamientoA(28) and (AlmacenamientoB(28) xor Carry27)) or (AlmacenamientoB(28) and Carry27); 

Resultado1(29) <= (AlmacenamientoA(29) and (AlmacenamientoB(29) xnor Carry28)) or (not AlmacenamientoA(29) and (AlmacenamientoB(29) xor Carry28)); 
Carry29 <= (AlmacenamientoA(29) and (AlmacenamientoB(29) xor Carry28)) or (AlmacenamientoB(29) and Carry28); 
 
Resultado1(30) <= (AlmacenamientoA(30) and (AlmacenamientoB(30) xnor Carry29)) or (not AlmacenamientoA(30) and (AlmacenamientoB(30) xor Carry29)); 
Carry30 <= (AlmacenamientoA(30) and (AlmacenamientoB(30) xor Carry29)) or (AlmacenamientoB(30) and Carry29); 

Resultado1(31) <= (AlmacenamientoA(31) and (AlmacenamientoB(31) xnor Carry30)) or (not AlmacenamientoA(31) and (AlmacenamientoB(31) xor Carry30)); 


-------SUBTRACT--------------

Complemento1(0) <= ((AlmacenamientoA(0) and (AlmacenamientoBN(0)xnor not AlmacI)) or (not AlmacenamientoA(0) and (AlmacenamientoBN(0) xor not AlmacI))); 
CarryZ0 <= (AlmacenamientoA(0) and (AlmacenamientoBN(0)));  

Complemento1(1) <= (AlmacenamientoA(1) and (AlmacenamientoBN(1) xnor CarryZ0)) or (not AlmacenamientoA(1) and (AlmacenamientoBN(1) xor CarryZ0)); 
CarryZ1 <= (AlmacenamientoA(1) and (AlmacenamientoBN(1) xor CarryZ0)) or (AlmacenamientoBN(1) and CarryZ0); 

Complemento1(2) <= (AlmacenamientoA(2)and (AlmacenamientoBN(2)xnor CarryZ1)) or (not AlmacenamientoA(2)and (AlmacenamientoBN(2)xor CarryZ1)); 
CarryZ2 <= (AlmacenamientoA(2)and (AlmacenamientoBN(2)xor CarryZ1)) or (AlmacenamientoBN(2)and CarryZ1); 

Complemento1(3) <= (AlmacenamientoA(3)and (AlmacenamientoBN(3)xnor CarryZ2)) or (not AlmacenamientoA(3)and  (AlmacenamientoBN(3)xor CarryZ2)); 
CarryZ3 <= (AlmacenamientoA(3)and (AlmacenamientoBN(3)xor CarryZ2)) or (AlmacenamientoBN(3)and CarryZ2); 

Complemento1(4) <= (AlmacenamientoA(4)and (AlmacenamientoBN(4)xnor CarryZ3)) or (not AlmacenamientoA(4)and (AlmacenamientoBN(4)xor CarryZ3)); 
CarryZ4 <= (AlmacenamientoA(4)and (AlmacenamientoBN(4)xor CarryZ3)) or (AlmacenamientoBN(4)and CarryZ3); 

Complemento1(5) <= (AlmacenamientoA(5) and (AlmacenamientoBN(5) xnor CarryZ4)) or (not AlmacenamientoA(5) and (AlmacenamientoBN(5) xor CarryZ4)); 
CarryZ5 <= (AlmacenamientoA(5) and (AlmacenamientoBN(5) xor CarryZ4)) or (AlmacenamientoBN(5) and CarryZ4); 

Complemento1(6) <= (AlmacenamientoA(6) and (AlmacenamientoBN(6) xnor CarryZ5)) or (not AlmacenamientoA(6) and (AlmacenamientoBN(6) xor CarryZ5)); 
CarryZ6 <= (AlmacenamientoA(6) and (AlmacenamientoBN(6) xor CarryZ5)) or (AlmacenamientoBN(6) and CarryZ5); 

Complemento1(7) <= (AlmacenamientoA(7) and (AlmacenamientoBN(7) xnor CarryZ6)) or (not AlmacenamientoA(7) and (AlmacenamientoBN(7) xor CarryZ6)); 
CarryZ7 <= (AlmacenamientoA(7) and (AlmacenamientoBN(7) xor CarryZ6)) or (AlmacenamientoBN(7) and CarryZ6); 

Complemento1(8) <= (AlmacenamientoA(8) and (AlmacenamientoBN(8) xnor CarryZ7)) or (not AlmacenamientoA(8) and (AlmacenamientoBN(8) xor CarryZ7)); 
CarryZ8 <= (AlmacenamientoA(8) and (AlmacenamientoBN(8) xor CarryZ7)) or (AlmacenamientoBN(8) and CarryZ7); 

Complemento1(9) <= (AlmacenamientoA(9) and (AlmacenamientoBN(9) xnor CarryZ8)) or (not AlmacenamientoA(9) and (AlmacenamientoBN(9) xor CarryZ8));
CarryZ9 <= (AlmacenamientoA(9) and (AlmacenamientoBN(9) xor CarryZ8)) or (AlmacenamientoBN(9) and CarryZ8); 

Complemento1(10) <= (AlmacenamientoA(10) and (AlmacenamientoBN(10) xnor CarryZ9)) or (not AlmacenamientoA(10) and (AlmacenamientoBN(10) xor CarryZ9)); 
CarryZ10 <= (AlmacenamientoA(10) and (AlmacenamientoBN(10) xor CarryZ9)) or (AlmacenamientoBN(10) and CarryZ9); 

Complemento1(11) <= (AlmacenamientoA(11) and (AlmacenamientoBN(11) xnor CarryZ10)) or (not AlmacenamientoA(11) and (AlmacenamientoBN(11) xor CarryZ10)); 
CarryZ11 <= (AlmacenamientoA(11) and (AlmacenamientoBN(11) xor CarryZ10)) or (AlmacenamientoBN(11) and CarryZ10); 

Complemento1(12) <= (AlmacenamientoA(12) and (AlmacenamientoBN(12) xnor CarryZ11)) or (not AlmacenamientoA(12) and (AlmacenamientoBN(12) xor CarryZ11)); 
CarryZ12 <= (AlmacenamientoA(12) and (AlmacenamientoBN(12) xor CarryZ11)) or (AlmacenamientoBN(12) and CarryZ11); 

Complemento1(13) <= (AlmacenamientoA(13) and (AlmacenamientoBN(13) xnor CarryZ12)) or (not AlmacenamientoA(13) and (AlmacenamientoBN(13) xor CarryZ12)); 
CarryZ13 <= (AlmacenamientoA(13) and (AlmacenamientoBN(13) xor CarryZ12)) or (AlmacenamientoBN(13) and CarryZ12); 

Complemento1(14) <= (AlmacenamientoA(14) and (AlmacenamientoBN(14) xnor CarryZ13)) or (not AlmacenamientoA(14) and (AlmacenamientoBN(14) xor CarryZ13)); 
CarryZ14 <= (AlmacenamientoA(14) and (AlmacenamientoBN(14) xor CarryZ13)) or (AlmacenamientoBN(14) and CarryZ13); 
 
Complemento1(15) <= (AlmacenamientoA(15) and (AlmacenamientoBN(15) xnor CarryZ14)) or (not AlmacenamientoA(15) and (AlmacenamientoBN(15) xor CarryZ14)); 
CarryZ15 <= (AlmacenamientoA(15) and (AlmacenamientoBN(15) xor CarryZ14)) or (AlmacenamientoBN(15) and CarryZ14); 

Complemento1(16) <= (AlmacenamientoA(16) and (AlmacenamientoBN(16) xnor CarryZ15)) or (not AlmacenamientoA(16) and (AlmacenamientoBN(16) xor CarryZ15)); 
CarryZ16 <= (AlmacenamientoA(16) and (AlmacenamientoBN(16) xor CarryZ15)) or (AlmacenamientoBN(16) and CarryZ15); 

Complemento1(17) <= (AlmacenamientoA(17)and (AlmacenamientoBN(17)xnor CarryZ16)) or (not AlmacenamientoA(17)and (AlmacenamientoBN(17)xor CarryZ16)); 
CarryZ17 <= (AlmacenamientoA(17)and (AlmacenamientoBN(17)xor CarryZ16)) or (AlmacenamientoBN(17)and CarryZ16); 

Complemento1(18) <= (AlmacenamientoA(18)and (AlmacenamientoBN(18)xnor CarryZ17)) or (not AlmacenamientoA(18)and  (AlmacenamientoBN(18)xor CarryZ17)); 
CarryZ18<= (AlmacenamientoA(18)and (AlmacenamientoBN(18)xor CarryZ17)) or (AlmacenamientoBN(18)and CarryZ17); 

Complemento1(19) <= (AlmacenamientoA(19)and (AlmacenamientoBN(19)xnor CarryZ18)) or (not AlmacenamientoA(19)and (AlmacenamientoBN(19)xor CarryZ18)); 
CarryZ19 <= (AlmacenamientoA(19)and (AlmacenamientoBN(19)xor CarryZ18)) or (AlmacenamientoBN(19)and CarryZ18); 

Complemento1(20) <= (AlmacenamientoA(20) and (AlmacenamientoBN(20) xnor CarryZ19)) or (not AlmacenamientoA(20) and (AlmacenamientoBN(20) xor CarryZ19)); 
CarryZ20 <= (AlmacenamientoA(20) and (AlmacenamientoBN(20) xor CarryZ19)) or (AlmacenamientoBN(20) and CarryZ19); 

Complemento1(21) <= (AlmacenamientoA(21) and (AlmacenamientoBN(21) xnor CarryZ20)) or (not AlmacenamientoA(21) and (AlmacenamientoBN(21) xor CarryZ20)); 
CarryZ21 <= (AlmacenamientoA(21) and (AlmacenamientoBN(21) xor CarryZ20)) or (AlmacenamientoBN(21) and CarryZ20); 

Complemento1(22) <= (AlmacenamientoA(22) and (AlmacenamientoBN(22) xnor CarryZ21)) or (not AlmacenamientoA(22) and (AlmacenamientoBN(22) xor CarryZ21)); 
CarryZ22 <= (AlmacenamientoA(22) and (AlmacenamientoBN(22) xor CarryZ21)) or (AlmacenamientoBN(22) and CarryZ21); 

Complemento1(23) <= (AlmacenamientoA(23) and (AlmacenamientoBN(23) xnor CarryZ22)) or (not AlmacenamientoA(23) and (AlmacenamientoBN(23) xor CarryZ22)); 
CarryZ23 <= (AlmacenamientoA(23) and (AlmacenamientoBN(23) xor CarryZ22)) or (AlmacenamientoBN(23) and CarryZ22); 
 
Complemento1(24) <= (AlmacenamientoA(24) and (AlmacenamientoBN(24) xnor CarryZ23)) or (not AlmacenamientoA(24) and (AlmacenamientoBN(24) xor CarryZ23)); 
CarryZ24 <= (AlmacenamientoA(24) and (AlmacenamientoBN(24) xor CarryZ23)) or (AlmacenamientoBN(24) and CarryZ23); 

Complemento1(25) <= (AlmacenamientoA(25) and (AlmacenamientoBN(25) xnor CarryZ24)) or (not AlmacenamientoA(25) and (AlmacenamientoBN(25) xor CarryZ24)); 
CarryZ25 <= (AlmacenamientoA(25) and (AlmacenamientoBN(25) xor CarryZ24)) or (AlmacenamientoBN(25) and CarryZ24); 

Complemento1(26) <= (AlmacenamientoA(26) and (AlmacenamientoBN(26) xnor CarryZ25)) or (not AlmacenamientoA(26) and (AlmacenamientoBN(26) xor CarryZ25)); 
CarryZ26 <= (AlmacenamientoA(26) and (AlmacenamientoBN(26) xor CarryZ25)) or (AlmacenamientoBN(26) and CarryZ25); 

Complemento1(27) <= (AlmacenamientoA(27) and (AlmacenamientoBN(27) xnor CarryZ26)) or (not AlmacenamientoA(27) and (AlmacenamientoBN(27) xor CarryZ26)); 
CarryZ27 <= (AlmacenamientoA(27) and (AlmacenamientoBN(27) xor CarryZ26)) or (AlmacenamientoBN(27) and CarryZ26); 

Complemento1(28) <= (AlmacenamientoA(28) and (AlmacenamientoBN(28) xnor CarryZ27)) or (not AlmacenamientoA(28) and (AlmacenamientoBN(28) xor CarryZ27)); 
CarryZ28 <= (AlmacenamientoA(28) and (AlmacenamientoBN(28) xor CarryZ27)) or (AlmacenamientoBN(28) and CarryZ27); 

Complemento1(29) <= (AlmacenamientoA(29) and (AlmacenamientoBN(29) xnor CarryZ28)) or (not AlmacenamientoA(29) and (AlmacenamientoBN(29) xor CarryZ28)); 
CarryZ29 <= (AlmacenamientoA(29) and (AlmacenamientoBN(29) xor CarryZ28)) or (AlmacenamientoBN(29) and CarryZ28); 
 
Complemento1(30) <= (AlmacenamientoA(30) and (AlmacenamientoBN(30) xnor CarryZ29)) or (not AlmacenamientoA(30) and (AlmacenamientoBN(30) xor CarryZ29)); 
CarryZ30 <= (AlmacenamientoA(30) and (AlmacenamientoBN(30) xor CarryZ29)) or (AlmacenamientoBN(30) and CarryZ29); 

Complemento1(31) <= (AlmacenamientoA(31) and (AlmacenamientoBN(31) xnor CarryZ30)) or (not AlmacenamientoA(31) and (AlmacenamientoBN(31) xor CarryZ30));






-----si carry es 1 se suma al primer bit sino se invierte el resultado---------------
Complemento2(0) <= ((Complemento1(0) and (Acarreo(0)xnor not AlmacI)) or (not Complemento1(0) and (Acarreo(0) xor not AlmacI))); 
CarryX0 <= (Complemento1(0) and (Acarreo(0)));  

Complemento2(1) <= (Complemento1(1) and (Acarreo(1) xnor CarryX0)) or (not Complemento1(1) and (Acarreo(1) xor CarryX0)); 
CarryX1 <= (Complemento1(1) and (Acarreo(1) xor CarryX0)) or (Acarreo(1) and CarryX0); 

Complemento2(2) <= (Complemento1(2)and (Acarreo(2)xnor CarryX1)) or (not Complemento1(2)and (Acarreo(2)xor CarryX1)); 
CarryX2 <= (Complemento1(2)and (Acarreo(2)xor CarryX1)) or (Acarreo(2)and CarryX1); 

Complemento2(3) <= (Complemento1(3)and (Acarreo(3)xnor CarryX2)) or (not Complemento1(3)and  (Acarreo(3)xor CarryX2)); 
CarryX3 <= (Complemento1(3)and (Acarreo(3)xor CarryX2)) or (Acarreo(3)and CarryX2); 

Complemento2(4) <= (Complemento1(4)and (Acarreo(4)xnor CarryX3)) or (not Complemento1(4)and (Acarreo(4)xor CarryX3)); 
CarryX4 <= (Complemento1(4)and (Acarreo(4)xor CarryX3)) or (Acarreo(4)and CarryX3); 

Complemento2(5) <= (Complemento1(5) and (Acarreo(5) xnor CarryX4)) or (not Complemento1(5) and (Acarreo(5) xor CarryX4)); 
CarryX5 <= (Complemento1(5) and (Acarreo(5) xor CarryX4)) or (Acarreo(5) and CarryX4); 

Complemento2(6) <= (Complemento1(6) and (Acarreo(6) xnor CarryX5)) or (not Complemento1(6) and (Acarreo(6) xor CarryX5)); 
CarryX6 <= (Complemento1(6) and (Acarreo(6) xor CarryX5)) or (Acarreo(6) and CarryX5); 

Complemento2(7) <= (Complemento1(7) and (Acarreo(7) xnor CarryX6)) or (not Complemento1(7) and (Acarreo(7) xor CarryX6)); 
CarryX7 <= (Complemento1(7) and (Acarreo(7) xor CarryX6)) or (Acarreo(7) and CarryX6); 

Complemento2(8) <= (Complemento1(8) and (Acarreo(8) xnor CarryX7)) or (not Complemento1(8) and (Acarreo(8) xor CarryX7)); 
CarryX8 <= (Complemento1(8) and (Acarreo(8) xor CarryX7)) or (Acarreo(8) and CarryX7); 

Complemento2(9) <= (Complemento1(9) and (Acarreo(9) xnor CarryX8)) or (not Complemento1(9) and (Acarreo(9) xor CarryX8));
CarryX9 <= (Complemento1(9) and (Acarreo(9) xor CarryX8)) or (Acarreo(9) and CarryX8); 

Complemento2(10) <= (Complemento1(10) and (Acarreo(10) xnor CarryX9)) or (not Complemento1(10) and (Acarreo(10) xor CarryX9)); 
CarryX10 <= (Complemento1(10) and (Acarreo(10) xor CarryX9)) or (Acarreo(10) and CarryX9); 

Complemento2(11) <= (Complemento1(11) and (Acarreo(11) xnor CarryX10)) or (not Complemento1(11) and (Acarreo(11) xor CarryX10)); 
CarryX11 <= (Complemento1(11) and (Acarreo(11) xor CarryX10)) or (Acarreo(11) and CarryX10); 

Complemento2(12) <= (Complemento1(12) and (Acarreo(12) xnor CarryX11)) or (not Complemento1(12) and (Acarreo(12) xor CarryX11)); 
CarryX12 <= (Complemento1(12) and (Acarreo(12) xor CarryX11)) or (Acarreo(12) and CarryX11); 

Complemento2(13) <= (Complemento1(13) and (Acarreo(13) xnor CarryX12)) or (not Complemento1(13) and (Acarreo(13) xor CarryX12)); 
CarryX13 <= (Complemento1(13) and (Acarreo(13) xor CarryX12)) or (Acarreo(13) and CarryX12); 

Complemento2(14) <= (Complemento1(14) and (Acarreo(14) xnor CarryX13)) or (not Complemento1(14) and (Acarreo(14) xor CarryX13)); 
CarryX14 <= (Complemento1(14) and (Acarreo(14) xor CarryX13)) or (Acarreo(14) and CarryX13); 
 
Complemento2(15) <= (Complemento1(15) and (Acarreo(15) xnor CarryX14)) or (not Complemento1(15) and (Acarreo(15) xor CarryX14)); 
CarryX15 <= (Complemento1(15) and (Acarreo(15) xor CarryX14)) or (Acarreo(15) and CarryX14); 

Complemento2(16) <= (Complemento1(16) and (Acarreo(16) xnor CarryX15)) or (not Complemento1(16) and (Acarreo(16) xor CarryX15)); 
CarryX16 <= (Complemento1(16) and (Acarreo(16) xor CarryX15)) or (Acarreo(16) and CarryX15); 

Complemento2(17) <= (Complemento1(17)and (Acarreo(17)xnor CarryX16)) or (not Complemento1(17)and (Acarreo(17)xor CarryX16)); 
CarryX17 <= (Complemento1(17)and (Acarreo(17)xor CarryX16)) or (Acarreo(17)and CarryX16); 

Complemento2(18) <= (Complemento1(18)and (Acarreo(18)xnor CarryX17)) or (not Complemento1(18)and  (Acarreo(18)xor CarryX17)); 
CarryX18<= (Complemento1(18)and (Acarreo(18)xor CarryX17)) or (Acarreo(18)and CarryX17); 

Complemento2(19) <= (Complemento1(19)and (Acarreo(19)xnor CarryX18)) or (not Complemento1(19)and (Acarreo(19)xor CarryX18)); 
CarryX19 <= (Complemento1(19)and (Acarreo(19)xor CarryX18)) or (Acarreo(19)and CarryX18); 

Complemento2(20) <= (Complemento1(20) and (Acarreo(20) xnor CarryX19)) or (not Complemento1(20) and (Acarreo(20) xor CarryX19)); 
CarryX20 <= (Complemento1(20) and (Acarreo(20) xor CarryX19)) or (Acarreo(20) and CarryX19); 

Complemento2(21) <= (Complemento1(21) and (Acarreo(21) xnor CarryX20)) or (not Complemento1(21) and (Acarreo(21) xor CarryX20)); 
CarryX21 <= (Complemento1(21) and (Acarreo(21) xor CarryX20)) or (Acarreo(21) and CarryX20); 

Complemento2(22) <= (Complemento1(22) and (Acarreo(22) xnor CarryX21)) or (not Complemento1(22) and (Acarreo(22) xor CarryX21)); 
CarryX22 <= (Complemento1(22) and (Acarreo(22) xor CarryX21)) or (Acarreo(22) and CarryX21); 

Complemento2(23) <= (Complemento1(23) and (Acarreo(23) xnor CarryX22)) or (not Complemento1(23) and (Acarreo(23) xor CarryX22)); 
CarryX23 <= (Complemento1(23) and (Acarreo(23) xor CarryX22)) or (Acarreo(23) and CarryX22); 
 
Complemento2(24) <= (Complemento1(24) and (Acarreo(24) xnor CarryX23)) or (not Complemento1(24) and (Acarreo(24) xor CarryX23)); 
CarryX24 <= (Complemento1(24) and (Acarreo(24) xor CarryX23)) or (Acarreo(24) and CarryX23); 

Complemento2(25) <= (Complemento1(25) and (Acarreo(25) xnor CarryX24)) or (not Complemento1(25) and (Acarreo(25) xor CarryX24)); 
CarryX25 <= (Complemento1(25) and (Acarreo(25) xor CarryX24)) or (Acarreo(25) and CarryX24); 

Complemento2(26) <= (Complemento1(26) and (Acarreo(26) xnor CarryX25)) or (not Complemento1(26) and (Acarreo(26) xor CarryX25)); 
CarryX26 <= (Complemento1(26) and (Acarreo(26) xor CarryX25)) or (Acarreo(26) and CarryX25); 

Complemento2(27) <= (Complemento1(27) and (Acarreo(27) xnor CarryX26)) or (not Complemento1(27) and (Acarreo(27) xor CarryX26)); 
CarryX27 <= (Complemento1(27) and (Acarreo(27) xor CarryX26)) or (Acarreo(27) and CarryX26); 

Complemento2(28) <= (Complemento1(28) and (Acarreo(28) xnor CarryX27)) or (not Complemento1(28) and (Acarreo(28) xor CarryX27)); 
CarryX28 <= (Complemento1(28) and (Acarreo(28) xor CarryX27)) or (Acarreo(28) and CarryX27); 

Complemento2(29) <= (Complemento1(29) and (Acarreo(29) xnor CarryX28)) or (not Complemento1(29) and (Acarreo(29) xor CarryX28)); 
CarryX29 <= (Complemento1(29) and (Acarreo(29) xor CarryX28)) or (Acarreo(29) and CarryX28); 
 
Complemento2(30) <= (Complemento1(30) and (Acarreo(30) xnor CarryX29)) or (not Complemento1(30) and (Acarreo(30) xor CarryX29)); 
CarryX30 <= (Complemento1(30) and (Acarreo(30) xor CarryX29)) or (Acarreo(30) and CarryX29); 

Complemento2(31) <= (Complemento1(31) and (Acarreo(31) xnor CarryX30)) or (not Complemento1(31) and (Acarreo(31) xor CarryX30));



resultado2(0)<=(CarryZ30 and complemento2(0)) or(not CarryZ30 and not complemento1(0));
resultado2(1)<=(CarryZ30 and complemento2(1)) or(not CarryZ30 and not complemento1(1));
resultado2(2)<=(CarryZ30 and complemento2(2)) or(not CarryZ30 and not complemento1(2));
resultado2(3)<=(CarryZ30 and complemento2(3)) or(not CarryZ30 and not complemento1(3));
resultado2(4)<=(CarryZ30 and complemento2(4)) or(not CarryZ30 and not complemento1(4));
resultado2(5)<=(CarryZ30 and complemento2(5)) or(not CarryZ30 and not complemento1(5));
resultado2(6)<=(CarryZ30 and complemento2(6)) or(not CarryZ30 and not complemento1(6));
resultado2(7)<=(CarryZ30 and complemento2(7)) or(not CarryZ30 and not complemento1(7));
resultado2(8)<=(CarryZ30 and complemento2(8)) or(not CarryZ30 and not complemento1(8));
resultado2(9)<=(CarryZ30 and complemento2(9)) or(not CarryZ30 and not complemento1(9));
resultado2(10)<=(CarryZ30 and complemento2(10)) or(not CarryZ30 and not complemento1(10));
resultado2(11)<=(CarryZ30 and complemento2(11)) or(not CarryZ30 and not complemento1(11));
resultado2(12)<=(CarryZ30 and complemento2(12)) or(not CarryZ30 and not complemento1(12));
resultado2(13)<=(CarryZ30 and complemento2(13)) or(not CarryZ30 and not complemento1(13));
resultado2(14)<=(CarryZ30 and complemento2(14)) or(not CarryZ30 and not complemento1(14));
resultado2(15)<=(CarryZ30 and complemento2(15)) or(not CarryZ30 and not complemento1(15));
resultado2(16)<=(CarryZ30 and complemento2(16)) or(not CarryZ30 and not complemento1(16));
resultado2(17)<=(CarryZ30 and complemento2(17)) or(not CarryZ30 and not complemento1(17));
resultado2(18)<=(CarryZ30 and complemento2(18)) or(not CarryZ30 and not complemento1(18));
resultado2(19)<=(CarryZ30 and complemento2(19)) or(not CarryZ30 and not complemento1(19));
resultado2(20)<=(CarryZ30 and complemento2(20)) or(not CarryZ30 and not complemento1(20));
resultado2(21)<=(CarryZ30 and complemento2(21)) or(not CarryZ30 and not complemento1(21));
resultado2(22)<=(CarryZ30 and complemento2(22)) or(not CarryZ30 and not complemento1(22));
resultado2(23)<=(CarryZ30 and complemento2(23)) or(not CarryZ30 and not complemento1(23));
resultado2(24)<=(CarryZ30 and complemento2(24)) or(not CarryZ30 and not complemento1(24));
resultado2(25)<=(CarryZ30 and complemento2(25)) or(not CarryZ30 and not complemento1(25));
resultado2(26)<=(CarryZ30 and complemento2(26)) or(not CarryZ30 and not complemento1(26));
resultado2(27)<=(CarryZ30 and complemento2(27)) or(not CarryZ30 and not complemento1(27));
resultado2(28)<=(CarryZ30 and complemento2(28)) or(not CarryZ30 and not complemento1(28));
resultado2(29)<=(CarryZ30 and complemento2(29)) or(not CarryZ30 and not complemento1(29));
resultado2(30)<=(CarryZ30 and complemento2(30)) or(not CarryZ30 and not complemento1(30));
resultado2(31)<=(CarryZ30 and complemento2(31)) or(not CarryZ30 and not complemento1(31));


-------AND------
Resultado3(0)   <= AlmacenamientoA(0) and AlmacenamientoB(0);    
Resultado3(1)   <= AlmacenamientoA(1) and AlmacenamientoB(1);    
Resultado3(2)   <= AlmacenamientoA(2) and AlmacenamientoB(2);    
Resultado3(3)   <= AlmacenamientoA(3) and AlmacenamientoB(3);    
Resultado3(4)   <= AlmacenamientoA(4) and AlmacenamientoB(4);    
Resultado3(5)   <= AlmacenamientoA(5) and AlmacenamientoB(5);    
Resultado3(6)   <= AlmacenamientoA(6) and AlmacenamientoB(6);    
Resultado3(7)   <= AlmacenamientoA(7) and AlmacenamientoB(7);    
Resultado3(8)   <= AlmacenamientoA(8) and AlmacenamientoB(8);    
Resultado3(9)   <= AlmacenamientoA(9) and AlmacenamientoB(9);    
Resultado3(10)  <= AlmacenamientoA(10) and AlmacenamientoB(10);    
Resultado3(11)  <= AlmacenamientoA(11) and AlmacenamientoB(11);    
Resultado3(12)  <= AlmacenamientoA(12) and AlmacenamientoB(12);    
Resultado3(13)  <= AlmacenamientoA(13) and AlmacenamientoB(13);    
Resultado3(14)  <= AlmacenamientoA(14) and AlmacenamientoB(14);    
Resultado3(15)  <= AlmacenamientoA(15) and AlmacenamientoB(15);    
Resultado3(16)  <= AlmacenamientoA(16) and AlmacenamientoB(16);    
Resultado3(17)  <= AlmacenamientoA(17) and AlmacenamientoB(17);   
Resultado3(18)  <= AlmacenamientoA(18) and AlmacenamientoB(18);    
Resultado3(19)  <= AlmacenamientoA(19) and AlmacenamientoB(19);    
Resultado3(20)  <= AlmacenamientoA(20) and AlmacenamientoB(20);    
Resultado3(21)  <= AlmacenamientoA(21) and AlmacenamientoB(21);    
Resultado3(22)  <= AlmacenamientoA(22) and AlmacenamientoB(22);    
Resultado3(23)  <= AlmacenamientoA(23) and AlmacenamientoB(23);    
Resultado3(24)  <= AlmacenamientoA(24) and AlmacenamientoB(24);    
Resultado3(25)  <= AlmacenamientoA(25) and AlmacenamientoB(25);    
Resultado3(26)  <= AlmacenamientoA(26) and AlmacenamientoB(26);    
Resultado3(27)  <= AlmacenamientoA(27) and AlmacenamientoB(27);    
Resultado3(28)  <= AlmacenamientoA(28) and AlmacenamientoB(28);    
Resultado3(29)  <= AlmacenamientoA(29) and AlmacenamientoB(29);    
Resultado3(30)  <= AlmacenamientoA(30) and AlmacenamientoB(30);    
Resultado3(31)  <= AlmacenamientoA(31) and AlmacenamientoB(31);

------OR---------
Resultado4(0)  <= AlmacenamientoA(0) or  AlmacenamientoB(0);    
Resultado4(1)  <= AlmacenamientoA(1) or AlmacenamientoB(1);    
Resultado4(2)  <= AlmacenamientoA(2) or AlmacenamientoB(2);    
Resultado4(3)  <= AlmacenamientoA(3) or AlmacenamientoB(3);    
Resultado4(4)  <= AlmacenamientoA(4) or AlmacenamientoB(4);    
Resultado4(5)  <= AlmacenamientoA(5) or AlmacenamientoB(5);    
Resultado4(6)  <= AlmacenamientoA(6) or AlmacenamientoB(6);    
Resultado4(7)  <= AlmacenamientoA(7) or AlmacenamientoB(7);    
Resultado4(8)  <= AlmacenamientoA(8) or AlmacenamientoB(8);    
Resultado4(9)  <= AlmacenamientoA(9) or AlmacenamientoB(9);    
Resultado4(10)  <= AlmacenamientoA(10) or AlmacenamientoB(10);    
Resultado4(11)  <= AlmacenamientoA(11) or AlmacenamientoB(11);    
Resultado4(12)  <= AlmacenamientoA(12) or AlmacenamientoB(12);    
Resultado4(13)  <= AlmacenamientoA(13) or AlmacenamientoB(13);    
Resultado4(14)  <= AlmacenamientoA(14) or AlmacenamientoB(14);    
Resultado4(15)  <= AlmacenamientoA(15) or AlmacenamientoB(15);    
Resultado4(16)  <= AlmacenamientoA(16) or AlmacenamientoB(16);    
Resultado4(17)  <= AlmacenamientoA(17) or AlmacenamientoB(17);   
Resultado4(18)  <= AlmacenamientoA(18) or AlmacenamientoB(18);    
Resultado4(19)  <= AlmacenamientoA(19) or AlmacenamientoB(19);    
Resultado4(20)  <= AlmacenamientoA(20) or AlmacenamientoB(20);    
Resultado4(21)  <= AlmacenamientoA(21) or AlmacenamientoB(21);    
Resultado4(22)  <= AlmacenamientoA(22) or AlmacenamientoB(22);    
Resultado4(23)  <= AlmacenamientoA(23) or AlmacenamientoB(23);    
Resultado4(24)  <= AlmacenamientoA(24) or AlmacenamientoB(24);    
Resultado4(25)  <= AlmacenamientoA(25) or AlmacenamientoB(25);    
Resultado4(26)  <= AlmacenamientoA(26) or AlmacenamientoB(26);    
Resultado4(27)  <= AlmacenamientoA(27) or AlmacenamientoB(27);    
Resultado4(28)  <= AlmacenamientoA(28) or AlmacenamientoB(28);    
Resultado4(29)  <= AlmacenamientoA(29) or AlmacenamientoB(29);    
Resultado4(30)  <= AlmacenamientoA(30) or AlmacenamientoB(30);    
Resultado4(31)  <= AlmacenamientoA(31) or AlmacenamientoB(31);

--------XOR---------
Resultado5(0)  <= AlmacenamientoA(0) xor  AlmacenamientoB(0);    
Resultado5(1)  <= AlmacenamientoA(1) xor AlmacenamientoB(1);    
Resultado5(2)  <= AlmacenamientoA(2) xor AlmacenamientoB(2);    
Resultado5(3)  <= AlmacenamientoA(3) xor AlmacenamientoB(3);    
Resultado5(4)  <= AlmacenamientoA(4) xor AlmacenamientoB(4);    
Resultado5(5)  <= AlmacenamientoA(5) xor AlmacenamientoB(5);    
Resultado5(6)  <= AlmacenamientoA(6) xor AlmacenamientoB(6);    
Resultado5(7)  <= AlmacenamientoA(7) xor AlmacenamientoB(7);    
Resultado5(8)  <= AlmacenamientoA(8) xor AlmacenamientoB(8);    
Resultado5(9)  <= AlmacenamientoA(9) xor AlmacenamientoB(9);    
Resultado5(10)  <= AlmacenamientoA(10) xor AlmacenamientoB(10);    
Resultado5(11)  <= AlmacenamientoA(11) xor AlmacenamientoB(11);    
Resultado5(12)  <= AlmacenamientoA(12) xor AlmacenamientoB(12);    
Resultado5(13)  <= AlmacenamientoA(13) xor AlmacenamientoB(13);    
Resultado5(14)  <= AlmacenamientoA(14) xor AlmacenamientoB(14);    
Resultado5(15)  <= AlmacenamientoA(15) xor AlmacenamientoB(15);    
Resultado5(16)  <= AlmacenamientoA(16) xor AlmacenamientoB(16);    
Resultado5(17)  <= AlmacenamientoA(17) xor AlmacenamientoB(17);   
Resultado5(18)  <= AlmacenamientoA(18) xor AlmacenamientoB(18);    
Resultado5(19)  <= AlmacenamientoA(19) xor AlmacenamientoB(19);    
Resultado5(20)  <= AlmacenamientoA(20) xor AlmacenamientoB(20);    
Resultado5(21)  <= AlmacenamientoA(21) xor AlmacenamientoB(21);    
Resultado5(22)  <= AlmacenamientoA(22) xor AlmacenamientoB(22);    
Resultado5(23)  <= AlmacenamientoA(23) xor AlmacenamientoB(23);    
Resultado5(24)  <= AlmacenamientoA(24) xor AlmacenamientoB(24);    
Resultado5(25)  <= AlmacenamientoA(25) xor AlmacenamientoB(25);    
Resultado5(26)  <= AlmacenamientoA(26) xor AlmacenamientoB(26);    
Resultado5(27)  <= AlmacenamientoA(27) xor AlmacenamientoB(27);    
Resultado5(28)  <= AlmacenamientoA(28) xor AlmacenamientoB(28);    
Resultado5(29)  <= AlmacenamientoA(29) xor AlmacenamientoB(29);    
Resultado5(30)  <= AlmacenamientoA(30) xor AlmacenamientoB(30);    
Resultado5(31)  <= AlmacenamientoA(31) xor AlmacenamientoB(31);


----------ROTATE R-----
Resultado6(0)<=(AlmacenamientoA(0) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(7) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(1)<=(AlmacenamientoA(1) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(8) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(2)<=(AlmacenamientoA(2) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(9) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(3)<=(AlmacenamientoA(3) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(10) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(4)<=(AlmacenamientoA(4) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(11) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(5)<=(AlmacenamientoA(5) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(12) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(6)<=(AlmacenamientoA(6) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(13) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(7)<=(AlmacenamientoA(7) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(14) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(8)<=(AlmacenamientoA(8) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(15) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(9)<=(AlmacenamientoA(9) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(16) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(10)<=(AlmacenamientoA(10) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(17) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(11)<=(AlmacenamientoA(11) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(18) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(12)<=(AlmacenamientoA(12) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(19) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(30)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(13)<=(AlmacenamientoA(13) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(20) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(31)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(14)<=(AlmacenamientoA(14) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(21) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(0)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(15)<=(AlmacenamientoA(15) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(22) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(1)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(16)<=(AlmacenamientoA(16) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(23) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(2)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(17)<=(AlmacenamientoA(17) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(24) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(3)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(18)<=(AlmacenamientoA(18) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(25) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(4)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(19)<=(AlmacenamientoA(19) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(26) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(5)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(20)<=(AlmacenamientoA(20) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(27) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(6)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(21)<=(AlmacenamientoA(21) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(28) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(7)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(22)<=(AlmacenamientoA(22) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(29) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(8)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(23)<=(AlmacenamientoA(23) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(30) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(9)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(24)<=(AlmacenamientoA(24) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(31) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(10)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(25)<=(AlmacenamientoA(25) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(0) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(11)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(26)<=(AlmacenamientoA(26) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(1) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(12)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(27)<=(AlmacenamientoA(27) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(0) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(13)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(28)<=(AlmacenamientoA(28) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(3) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(14)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(29)<=(AlmacenamientoA(29) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(30)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(4) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(15)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(30)<=(AlmacenamientoA(30) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(31)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(5) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(6)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(15)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(16)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(17)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(27)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(28)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(29)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
Resultado6(31)<=(AlmacenamientoA(31) AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(0)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(1)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(2)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(3)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(4)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR ( AlmacenamientoA(6) AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(7)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(8)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(9)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(10)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(11)AND (not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(12)AND (AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(13)AND (not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(14)AND (AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(16)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR  (AlmacenamientoA(17)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(18)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(19)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(20)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(21)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(22)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND not AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(23)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(24)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(25)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(26)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND not AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(27)AND(not AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR  (AlmacenamientoA(28)AND(AlmacenamientoB(0) AND not AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4))) OR (AlmacenamientoA(29)AND(not AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)))OR (AlmacenamientoA(30)AND(AlmacenamientoB(0) AND AlmacenamientoB(1)AND AlmacenamientoB(2) AND AlmacenamientoB(3) AND AlmacenamientoB(4)));
----------END--ROTATE R------


-----SHIFT R-------- 
Resultado7(0)<=(AlmacenamientoA(0)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(1) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(2) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(3) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(7)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(18) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(1)<=(AlmacenamientoA(1)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(2) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(3) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(8)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(19) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0) AND (AlmacenamientoB(1)  AND  AlmacenamientoB(2) AND  AlmacenamientoB(3)   AND  AlmacenamientoB(4))));
Resultado7(2)<=(AlmacenamientoA(2)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(3) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(9)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(20) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(3)<=(AlmacenamientoA(3)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(4) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(10)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(21) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(4)<=(AlmacenamientoA(4)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(5) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(11)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(22) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(5)<=(AlmacenamientoA(5)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(6) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(12)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(23) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(6)<=(AlmacenamientoA(6)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(7) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(13)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(24) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(7)<=(AlmacenamientoA(7)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(8) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(14)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(25) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(8)<=(AlmacenamientoA(8)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(9) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(15)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(26) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(9)<=(AlmacenamientoA(9)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(10) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(16)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(27) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(10)<=(AlmacenamientoA(10)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(17)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(28) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(11)<=(AlmacenamientoA(11)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(12) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(18)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(29) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(12)<=(AlmacenamientoA(12)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(19)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(30) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(13)<=(AlmacenamientoA(13)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(20)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(14)<=(AlmacenamientoA(14)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(15) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(21)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(15)<=(AlmacenamientoA(15)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(16) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(22)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(16)<=(AlmacenamientoA(16)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(17) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(23)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(17)<=(AlmacenamientoA(17)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(18) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(24)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(18)<=(AlmacenamientoA(18)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(19) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(25)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(19)<=(AlmacenamientoA(19)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(20) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(26)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(20)<=(AlmacenamientoA(20)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(21) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(27)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(21)<=(AlmacenamientoA(21)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(22) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(28)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(22)<=(AlmacenamientoA(22)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(23) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(29)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(23)<=(AlmacenamientoA(23)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(24) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(30)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(24)<=(AlmacenamientoA(24)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(25) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(25)<=(AlmacenamientoA(25)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(26) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(26)<=(AlmacenamientoA(26)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(27) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(27)<=(AlmacenamientoA(27)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(28) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(28)<=(AlmacenamientoA(28)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(29) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(29)<=(AlmacenamientoA(29)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(30) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(30)<=(AlmacenamientoA(30)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(11) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(13) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(14)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
Resultado7(31)<=(AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR ( AlmacenamientoA(31)  AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND  (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  not AlmacenamientoB(4))) OR (AlmacenamientoA(31)  AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR  (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  not AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  not AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)))OR  (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  not AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4))) OR (AlmacenamientoA(31) AND (not AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)) )OR (AlmacenamientoA(31) AND (AlmacenamientoB(0)  AND  AlmacenamientoB(1) AND  AlmacenamientoB(2)  AND  AlmacenamientoB(3)  AND  AlmacenamientoB(4)));
-----END--SHIFT R--------




---------HABILTAR_SALIDA DE ALU-------------------------------------------------------
OpcodeSuma<=(not ALU_Control(0) and not ALU_Control(1) and not ALU_Control(2));--000---
OpcodeResta<=(ALU_Control(0) and not ALU_Control(1) and not ALU_Control(2));--100--
OpcodeAnd<=(not ALU_Control(0) and  ALU_Control(1) and not ALU_Control(2));--010--
OpcodeOr<=( ALU_Control(0) and  ALU_Control(1) and not ALU_Control(2));--110--
OpcodeXor<=(not ALU_Control(0) and not ALU_Control(1) and  ALU_Control(2));--001--
OpcodeRotate<=(ALU_Control(0) and not ALU_Control(1) and  ALU_Control(2));--101--
OpcodeShift<=(not ALU_Control(0) and  ALU_Control(1) and  ALU_Control(2));--011--
--------------------------------------------------------------------------------------
Salida1(0)  <= Resultado1(0) and  OpcodeSuma;    
Salida1(1)  <= Resultado1(1) and OpcodeSuma;    
Salida1(2)  <= Resultado1(2) and OpcodeSuma;    
Salida1(3)  <= Resultado1(3) and OpcodeSuma;    
Salida1(4)  <= Resultado1(4) and OpcodeSuma;    
Salida1(5)  <= Resultado1(5) and OpcodeSuma;    
Salida1(6)  <= Resultado1(6) and OpcodeSuma;    
Salida1(7)  <= Resultado1(7) and OpcodeSuma;    
Salida1(8)  <= Resultado1(8) and OpcodeSuma;    
Salida1(9)  <= Resultado1(9) and OpcodeSuma;    
Salida1(10)  <= Resultado1(10) and OpcodeSuma;    
Salida1(11)  <= Resultado1(11) and OpcodeSuma;    
Salida1(12)  <= Resultado1(12) and OpcodeSuma;    
Salida1(13)  <= Resultado1(13) and OpcodeSuma;    
Salida1(14)  <= Resultado1(14) and OpcodeSuma;    
Salida1(15)  <= Resultado1(15) and OpcodeSuma;    
Salida1(16)  <= Resultado1(16) and OpcodeSuma;    
Salida1(17)  <= Resultado1(17) and OpcodeSuma;   
Salida1(18)  <= Resultado1(18) and OpcodeSuma;    
Salida1(19)  <= Resultado1(19) and OpcodeSuma;    
Salida1(20)  <= Resultado1(20) and OpcodeSuma;    
Salida1(21)  <= Resultado1(21) and OpcodeSuma;    
Salida1(22)  <= Resultado1(22) and OpcodeSuma;    
Salida1(23)  <= Resultado1(23) and OpcodeSuma;    
Salida1(24)  <= Resultado1(24) and OpcodeSuma;    
Salida1(25)  <= Resultado1(25) and OpcodeSuma;    
Salida1(26)  <= Resultado1(26) and OpcodeSuma;    
Salida1(27)  <= Resultado1(27) and OpcodeSuma;    
Salida1(28)  <= Resultado1(28) and OpcodeSuma;    
Salida1(29)  <= Resultado1(29) and OpcodeSuma;    
Salida1(30)  <= Resultado1(30) and OpcodeSuma;    
Salida1(31)  <= Resultado1(31) and OpcodeSuma;

Salida2(0)  <= Resultado2(0) and  OpcodeResta;    
Salida2(1)  <= Resultado2(1) and OpcodeResta;    
Salida2(2)  <= Resultado2(2) and OpcodeResta;    
Salida2(3)  <= Resultado2(3) and OpcodeResta;    
Salida2(4)  <= Resultado2(4) and OpcodeResta;    
Salida2(5)  <= Resultado2(5) and OpcodeResta;    
Salida2(6)  <= Resultado2(6) and OpcodeResta;    
Salida2(7)  <= Resultado2(7) and OpcodeResta;    
Salida2(8)  <= Resultado2(8) and OpcodeResta;    
Salida2(9)  <= Resultado2(9) and OpcodeResta;    
Salida2(10)  <= Resultado2(10) and OpcodeResta;    
Salida2(11)  <= Resultado2(11) and OpcodeResta;    
Salida2(12)  <= Resultado2(12) and OpcodeResta;    
Salida2(13)  <= Resultado2(13) and OpcodeResta;    
Salida2(14)  <= Resultado2(14) and OpcodeResta;    
Salida2(15)  <= Resultado2(15) and OpcodeResta;    
Salida2(16)  <= Resultado2(16) and OpcodeResta;    
Salida2(17)  <= Resultado2(17) and OpcodeResta;   
Salida2(18)  <= Resultado2(18) and OpcodeResta;    
Salida2(19)  <= Resultado2(19) and OpcodeResta;    
Salida2(20)  <= Resultado2(20) and OpcodeResta;    
Salida2(21)  <= Resultado2(21) and OpcodeResta;    
Salida2(22)  <= Resultado2(22) and OpcodeResta;    
Salida2(23)  <= Resultado2(23) and OpcodeResta;    
Salida2(24)  <= Resultado2(24) and OpcodeResta;    
Salida2(25)  <= Resultado2(25) and OpcodeResta;    
Salida2(26)  <= Resultado2(26) and OpcodeResta;    
Salida2(27)  <= Resultado2(27) and OpcodeResta;    
Salida2(28)  <= Resultado2(28) and OpcodeResta;    
Salida2(29)  <= Resultado2(29) and OpcodeResta;    
Salida2(30)  <= Resultado2(30) and OpcodeResta;    
Salida2(31)  <= Resultado2(31) and OpcodeResta;


Salida3(0)  <= Resultado3(0) and  OpcodeAnd;    
Salida3(1)  <= Resultado3(1) and OpcodeAnd;    
Salida3(2)  <= Resultado3(2) and OpcodeAnd;    
Salida3(3)  <= Resultado3(3) and OpcodeAnd;    
Salida3(4)  <= Resultado3(4) and OpcodeAnd;    
Salida3(5)  <= Resultado3(5) and OpcodeAnd;    
Salida3(6)  <= Resultado3(6) and OpcodeAnd;    
Salida3(7)  <= Resultado3(7) and OpcodeAnd;    
Salida3(8)  <= Resultado3(8) and OpcodeAnd;    
Salida3(9)  <= Resultado3(9) and OpcodeAnd;    
Salida3(10)  <= Resultado3(10) and OpcodeAnd;    
Salida3(11)  <= Resultado3(11) and OpcodeAnd;    
Salida3(12)  <= Resultado3(12) and OpcodeAnd;    
Salida3(13)  <= Resultado3(13) and OpcodeAnd;    
Salida3(14)  <= Resultado3(14) and OpcodeAnd;    
Salida3(15)  <= Resultado3(15) and OpcodeAnd;    
Salida3(16)  <= Resultado3(16) and OpcodeAnd;    
Salida3(17)  <= Resultado3(17) and OpcodeAnd;   
Salida3(18)  <= Resultado3(18) and OpcodeAnd;    
Salida3(19)  <= Resultado3(19) and OpcodeAnd;    
Salida3(20)  <= Resultado3(20) and OpcodeAnd;    
Salida3(21)  <= Resultado3(21) and OpcodeAnd;    
Salida3(22)  <= Resultado3(22) and OpcodeAnd;    
Salida3(23)  <= Resultado3(23) and OpcodeAnd;    
Salida3(24)  <= Resultado3(24) and OpcodeAnd;    
Salida3(25)  <= Resultado3(25) and OpcodeAnd;    
Salida3(26)  <= Resultado3(26) and OpcodeAnd;    
Salida3(27)  <= Resultado3(27) and OpcodeAnd;    
Salida3(28)  <= Resultado3(28) and OpcodeAnd;    
Salida3(29)  <= Resultado3(29) and OpcodeAnd;    
Salida3(30)  <= Resultado3(30) and OpcodeAnd;    
Salida3(31)  <= Resultado3(31) and OpcodeAnd;


Salida4(0)  <= Resultado4(0) and  OpcodeOr;    
Salida4(1)  <= Resultado4(1) and OpcodeOr;    
Salida4(2)  <= Resultado4(2) and OpcodeOr;    
Salida4(3)  <= Resultado4(3) and OpcodeOr;    
Salida4(4)  <= Resultado4(4) and OpcodeOr;    
Salida4(5)  <= Resultado4(5) and OpcodeOr;    
Salida4(6)  <= Resultado4(6) and OpcodeOr;    
Salida4(7)  <= Resultado4(7) and OpcodeOr;    
Salida4(8)  <= Resultado4(8) and OpcodeOr;    
Salida4(9)  <= Resultado4(9) and OpcodeOr;    
Salida4(10)  <= Resultado4(10) and OpcodeOr;    
Salida4(11)  <= Resultado4(11) and OpcodeOr;    
Salida4(12)  <= Resultado4(12) and OpcodeOr;    
Salida4(13)  <= Resultado4(13) and OpcodeOr;    
Salida4(14)  <= Resultado4(14) and OpcodeOr;    
Salida4(15)  <= Resultado4(15) and OpcodeOr;    
Salida4(16)  <= Resultado4(16) and OpcodeOr;    
Salida4(17)  <= Resultado4(17) and OpcodeOr;   
Salida4(18)  <= Resultado4(18) and OpcodeOr;    
Salida4(19)  <= Resultado4(19) and OpcodeOr;    
Salida4(20)  <= Resultado4(20) and OpcodeOr;    
Salida4(21)  <= Resultado4(21) and OpcodeOr;    
Salida4(22)  <= Resultado4(22) and OpcodeOr;    
Salida4(23)  <= Resultado4(23) and OpcodeOr;    
Salida4(24)  <= Resultado4(24) and OpcodeOr;    
Salida4(25)  <= Resultado4(25) and OpcodeOr;    
Salida4(26)  <= Resultado4(26) and OpcodeOr;    
Salida4(27)  <= Resultado4(27) and OpcodeOr;    
Salida4(28)  <= Resultado4(28) and OpcodeOr;    
Salida4(29)  <= Resultado4(29) and OpcodeOr;    
Salida4(30)  <= Resultado4(30) and OpcodeOr;    
Salida4(31)  <= Resultado4(31) and OpcodeOr;


Salida5(0)  <= Resultado5(0) and  OpcodeXor;    
Salida5(1)  <= Resultado5(1) and OpcodeXor;    
Salida5(2)  <= Resultado5(2) and OpcodeXor;    
Salida5(3)  <= Resultado5(3) and OpcodeXor;    
Salida5(4)  <= Resultado5(4) and OpcodeXor;    
Salida5(5)  <= Resultado5(5) and OpcodeXor;    
Salida5(6)  <= Resultado5(6) and OpcodeXor;    
Salida5(7)  <= Resultado5(7) and OpcodeXor;    
Salida5(8)  <= Resultado5(8) and OpcodeXor;    
Salida5(9)  <= Resultado5(9) and OpcodeXor;    
Salida5(10)  <= Resultado5(10) and OpcodeXor;    
Salida5(11)  <= Resultado5(11) and OpcodeXor;    
Salida5(12)  <= Resultado5(12) and OpcodeXor;    
Salida5(13)  <= Resultado5(13) and OpcodeXor;    
Salida5(14)  <= Resultado5(14) and OpcodeXor;    
Salida5(15)  <= Resultado5(15) and OpcodeXor;    
Salida5(16)  <= Resultado5(16) and OpcodeXor;    
Salida5(17)  <= Resultado5(17) and OpcodeXor;   
Salida5(18)  <= Resultado5(18) and OpcodeXor;    
Salida5(19)  <= Resultado5(19) and OpcodeXor;    
Salida5(20)  <= Resultado5(20) and OpcodeXor;    
Salida5(21)  <= Resultado5(21) and OpcodeXor;    
Salida5(22)  <= Resultado5(22) and OpcodeXor;    
Salida5(23)  <= Resultado5(23) and OpcodeXor;    
Salida5(24)  <= Resultado5(24) and OpcodeXor;    
Salida5(25)  <= Resultado5(25) and OpcodeXor;    
Salida5(26)  <= Resultado5(26) and OpcodeXor;    
Salida5(27)  <= Resultado5(27) and OpcodeXor;    
Salida5(28)  <= Resultado5(28) and OpcodeXor;    
Salida5(29)  <= Resultado5(29) and OpcodeXor;    
Salida5(30)  <= Resultado5(30) and OpcodeXor;    
Salida5(31)  <= Resultado5(31) and OpcodeXor;


Salida6(0)  <= Resultado6(0) and  OpcodeRotate;    
Salida6(1)  <= Resultado6(1) and OpcodeRotate;    
Salida6(2)  <= Resultado6(2) and OpcodeRotate;    
Salida6(3)  <= Resultado6(3) and OpcodeRotate;    
Salida6(4)  <= Resultado6(4) and OpcodeRotate;    
Salida6(5)  <= Resultado6(5) and OpcodeRotate;    
Salida6(6)  <= Resultado6(6) and OpcodeRotate;    
Salida6(7)  <= Resultado6(7) and OpcodeRotate;    
Salida6(8)  <= Resultado6(8) and OpcodeRotate;    
Salida6(9)  <= Resultado6(9) and OpcodeRotate;    
Salida6(10)  <= Resultado6(10) and OpcodeRotate;    
Salida6(11)  <= Resultado6(11) and OpcodeRotate;    
Salida6(12)  <= Resultado6(12) and OpcodeRotate;    
Salida6(13)  <= Resultado6(13) and OpcodeRotate;    
Salida6(14)  <= Resultado6(14) and OpcodeRotate;    
Salida6(15)  <= Resultado6(15) and OpcodeRotate;    
Salida6(16)  <= Resultado6(16) and OpcodeRotate;    
Salida6(17)  <= Resultado6(17) and OpcodeRotate;   
Salida6(18)  <= Resultado6(18) and OpcodeRotate;    
Salida6(19)  <= Resultado6(19) and OpcodeRotate;    
Salida6(20)  <= Resultado6(20) and OpcodeRotate;    
Salida6(21)  <= Resultado6(21) and OpcodeRotate;    
Salida6(22)  <= Resultado6(22) and OpcodeRotate;    
Salida6(23)  <= Resultado6(23) and OpcodeRotate;    
Salida6(24)  <= Resultado6(24) and OpcodeRotate;    
Salida6(25)  <= Resultado6(25) and OpcodeRotate;    
Salida6(26)  <= Resultado6(26) and OpcodeRotate;    
Salida6(27)  <= Resultado6(27) and OpcodeRotate;    
Salida6(28)  <= Resultado6(28) and OpcodeRotate;    
Salida6(29)  <= Resultado6(29) and OpcodeRotate;    
Salida6(30)  <= Resultado6(30) and OpcodeRotate;    
Salida6(31)  <= Resultado6(31) and OpcodeRotate;

Salida7(0)  <= Resultado7(0) and  OpcodeShift;    
Salida7(1)  <= Resultado7(1) and OpcodeShift;    
Salida7(2)  <= Resultado7(2) and OpcodeShift;    
Salida7(3)  <= Resultado7(3) and OpcodeShift;    
Salida7(4)  <= Resultado7(4) and OpcodeShift;    
Salida7(5)  <= Resultado7(5) and OpcodeShift;    
Salida7(6)  <= Resultado7(6) and OpcodeShift;    
Salida7(7)  <= Resultado7(7) and OpcodeShift;    
Salida7(8)  <= Resultado7(8) and OpcodeShift;    
Salida7(9)  <= Resultado7(9) and OpcodeShift;    
Salida7(10)  <= Resultado7(10) and OpcodeShift;    
Salida7(11)  <= Resultado7(11) and OpcodeShift;    
Salida7(12)  <= Resultado7(12) and OpcodeShift;    
Salida7(13)  <= Resultado7(13) and OpcodeShift;    
Salida7(14)  <= Resultado7(14) and OpcodeShift;    
Salida7(15)  <= Resultado7(15) and OpcodeShift;    
Salida7(16)  <= Resultado7(16) and OpcodeShift;    
Salida7(17)  <= Resultado7(17) and OpcodeShift;   
Salida7(18)  <= Resultado7(18) and OpcodeShift;    
Salida7(19)  <= Resultado7(19) and OpcodeShift;    
Salida7(20)  <= Resultado7(20) and OpcodeShift;    
Salida7(21)  <= Resultado7(21) and OpcodeShift;    
Salida7(22)  <= Resultado7(22) and OpcodeShift;    
Salida7(23)  <= Resultado7(23) and OpcodeShift;    
Salida7(24)  <= Resultado7(24) and OpcodeShift;    
Salida7(25)  <= Resultado7(25) and OpcodeShift;    
Salida7(26)  <= Resultado7(26) and OpcodeShift;    
Salida7(27)  <= Resultado7(27) and OpcodeShift;    
Salida7(28)  <= Resultado7(28) and OpcodeShift;    
Salida7(29)  <= Resultado7(29) and OpcodeShift;    
Salida7(30)  <= Resultado7(30) and OpcodeShift;    
Salida7(31)  <= Resultado7(31) and OpcodeShift;
----------------------Salidas de ALU32---------------------------------------------------------
Equal_Than<=not Resultado2(0) and not Resultado2(1) and not Resultado2(2) and not Resultado2(3) and not Resultado2(4) and not Resultado2(5) and not Resultado2(6) and not Resultado2(7) and not Resultado2(8) and not Resultado2(9) and not Resultado2(10) and not Resultado2(11) and not Resultado2(12) and not Resultado2(13) and not Resultado2(14) and not Resultado2(15) and not Resultado2(16) and not Resultado2(17) and not Resultado2(18) and not Resultado2(19) and not Resultado2(20) and not Resultado2(21) and not Resultado2(22) and not Resultado2(23) and not Resultado2(24) and not Resultado2(25) and not Resultado2(26) and not Resultado2(27) and not Resultado2(28) and not Resultado2(29) and not Resultado2(30) and not Resultado2(31);
Larger_Than<=not ((AlmacenamientoA(31) XOR complemento2(31)) or (AlmacenamientoA(31) XOR complemento1(31)));
Less_Than<=not Larger_Than;
Not_Equal_Than<=not Equal_Than; 
SALIDA_ALU2<=(Equal_Than AND (ALU_Control2(0) and not ALU_Control2(1) and not ALU_Control2(2)and not ALU_Control2(3)))OR(Larger_Than AND (not ALU_Control2(0) and ALU_Control2(1) and not ALU_Control2(2)and not ALU_Control2(3)))OR(Less_Than AND (not ALU_Control2(0) and not ALU_Control2(1) and ALU_Control2(2)and not ALU_Control2(3))) or (Not_Equal_Than AND (not ALU_Control2(0) and not ALU_Control2(1) and not ALU_Control2(2) and  ALU_Control2(3)));
Salida_ALU1<=Salida1 or Salida2 or Salida3 or Salida4 or Salida5 or Salida6 or Salida7;
---prueba---
--igual<=Equal_Than;
--mayor<=Larger_Than;
--menor<=Less_Than;
---noigual<=Not_Equal_Than;
--restasalida<=Resultado2;
--twocomple<=complemento2;
--onecomple<=complemento1;
----------------
end ALU32Arch;

