--PONTIFICIA_UNIVERSIDAD_JAVERIANA-- 
--VHDL DE ROM-- 
--DISEÑADOR: DANIEL_FAJARDO-- 
--6/10/2020--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity ROM is
    generic(
        G_width     :integer := 15;
        G_word_size :integer := 32;
        G_length    :integer := 10
    );
    port(
        clk: in std_logic;
        addr: in std_logic_vector(G_width - 1 downto 0);
        dout: out std_logic_vector(G_word_size- 1 downto 0)
    ); 
end ROM;

architecture Behavioral of ROM is
    type rom_type is array (0 to 32767) of std_logic_vector(G_word_size- 1  downto 0);
    signal ROM: rom_type := (
        0      => "00000000000000000000000000000011", --1L
        1      => "00000000000000000001000010000011", --2L
        2      => "00000000000000000010000100000011", --3L
        3      => "00000000000000000011000110000011", --4L
        4      => "00000000000000000100001000000011", --5L
        5      => "00000000000000000101001010000011", --6L
        6      => "00000000000000000110001100000011", --7L
        7      => "00000000000000000111001110000011", --8L
        8      => "00000000000000000000101100000011", --9L
        9      => "00000000000000000000101100000011", --L
        10     => "00000000000000000000101100000011",
        11     => "00000000000011111000101100000011",
        12     => "00000000000011111000101100000011",
        13     => "00000000000011111000101100000011",
        14     => "00000000000011111000101100000011",
        15     => "00000000000011111000101100000011",
        16     => "00000000000011111000101100000011",
        17     => "00000001010110110101001001100011", --B
        18     => "00000000000000000000000000000011", --lL
        19     => "00000000000000000001000010000011", --1
        20     => "00000000000000000010000100000011", --2
        21     => "00000000000000000011000110000011", --3
        22     => "00000000000000000100001000000011", --4
        23     => "00000000000000000101001010000011", --5
        24     => "00000000000000000110001100000011", --7
        25     => "00000000100000000000111010010011", --I
        26     => "00000000000000000000000000000011", --L
        27     => "00000000000000000001000010000011", --L2--
        28     => "00000000001000000000101100000011",
        29     => "00000000001111110000101010000011",
        30     => "00000000010000000000101100000011",
        31     => "00000000010100000000101010000011",
        32     => "00000000011000000000101100000011",
        33     => "00000000011100000000101010000011",
        34     => "00000000100000000000101010000011",
        35     => "00000000100100000000101100000011",
        36     => "00000000101000000000101010000011",
        37     => "00000000101000000000101010000011",
        38     => "00000000101100000000101010000011",
        39     => "00000000110000000000101010000011",
        40     => "00000000000000000000111111111111", --sw
        41     => "00000000111000000000101010000011",
        42     => "00000000111100000000101010000011",
        others => "00000000000000000000000000110011"  --R
    );
begin
    process (clk)
    begin
        if rising_edge(clk) then
            dout <= ROM(to_integer(unsigned(addr(G_length - 1 downto 0))));
        end if;
    end process;
end Behavioral;
